module map(addr, data);
    input  [3:0] addr;  // addr = {coll, idx}
    output reg [7:0] data; // 輸出的綠燈資料 (1=牆壁/亮, 0=路徑/暗)

    always@(addr) begin
        case(addr)
            // ==========================================
            // Part 1: 正常遊戲模式 (coll=0, addr=0~7)
            // 這裡定義迷宮的牆壁。 "1" 代表牆壁 (綠燈亮)，"0" 代表路 (暗)
            // ==========================================
            4'd0 : data = 8'b1111_1111; // 第 0 列: 上方牆壁
            4'd1 : data = 8'b1000_0001; // 第 1 列: 左右有牆，中間是路
            4'd2 : data = 8'b1000_0001; // 第 2 列
            4'd3 : data = 8'b1001_1001; // 第 3 列: 中間加一些障礙物
            4'd4 : data = 8'b1000_0001; // 第 4 列
            4'd5 : data = 8'b1000_0001; // 第 5 列
            4'd6 : data = 8'b1000_0001; // 第 6 列
            4'd7 : data = 8'b1111_0001; // 第 7 列: 下方牆壁 (留一個出口在 bit 1~3)

            // ==========================================
            // Part 2: 碰撞模式 (coll=1, addr=8~15)
            // 當發生碰撞時，addr 會加上 8 (bit 3 變 1)
            // 根據 PPT ，撞到時全亮
            // ==========================================
            4'd8 : data = 8'b1111_1111;
            4'd9 : data = 8'b1111_1111;
            4'd10: data = 8'b1111_1111;
            4'd11: data = 8'b1111_1111;
            4'd12: data = 8'b1111_1111;
            4'd13: data = 8'b1111_1111;
            4'd14: data = 8'b1111_1111;
            4'd15: data = 8'b1111_1111;

            default: data = 8'b0000_0000;
        endcase
    end
endmodule